netcdf filter_input_saw {
dimensions:
	member = 80 ;
	metadatalength = 32 ;
	location = 10 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double concentration(time, member, location) ;
		concentration:long_name = "tracer concentration" ;
		concentration:units = "mass" ;

	double mean_source(time, member, location) ;
		mean_source:long_name = "mean source" ;
		mean_source:units = "mass/timestep" ;

	double source(time, member, location) ;
		source:long_name = "source" ;
		source:units = "mass/timestep" ;

	double source_phase(time, member, location) ;
		source_phase:long_name = "source phase" ;
		source_phase:units = "radians" ;

	double wind(time, member, location) ;
		wind:long_name = "wind" ;
		wind:units = "gridpoints/timestep" ;

	double concentration_priorinf_mean(time, location) ;
		concentration_priorinf_mean:long_name = "prior inflation value for concentration" ;

	double mean_source_priorinf_mean(time, location) ;
		mean_source_priorinf_mean:long_name = "prior inflation value for mean source" ;

	double source_phase_priorinf_mean(time, location) ;
		source_phase_priorinf_mean:long_name = "prior inflation value for source phase" ;

	double source_priorinf_mean(time, location) ;
		source_priorinf_mean:long_name = "prior inflation value for source" ;

	double wind_priorinf_mean(time, location) ;
		wind_priorinf_mean:long_name = "prior inflation value for wind" ;

	double concentration_priorinf_sd(time, location) ;
		concentration_priorinf_sd:long_name = "prior inflation standard deviation for concentration" ;

	double mean_source_priorinf_sd(time, location) ;
		mean_source_priorinf_sd:long_name = "prior inflation standard deviation for mean source" ;

	double source_phase_priorinf_sd(time, location) ;
		source_phase_priorinf_sd:long_name = "prior inflation standard deviation for source phase" ;

	double source_priorinf_sd(time, location) ;
		source_priorinf_sd:long_name = "prior inflation standard deviation for source" ;

	double wind_priorinf_sd(time, location) ;
		wind_priorinf_sd:long_name = "prior inflation standard deviation for wind" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;
		location:axis = "X" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

	double advance_to_time ;
		advance_to_time:long_name = "desired time at end of the next model advance" ;
		advance_to_time:axis = "T" ;
		advance_to_time:cartesian_axis = "T" ;
		advance_to_time:calendar = "none" ;
		advance_to_time:units = "days" ;

// global attributes:
		:title = "an ensemble of spun-up model states" ;
                :version = "$Id: filter_input_saw.cdl 11441 2017-04-06 22:00:44Z nancy@ucar.edu $" ;
                :description = "Saw tooth pattern for mean source at grid points 1 3 and 5" ;
		:model = "simple_advection" ;
		:destruction_rate = 5.555556e-05 ;
		:history = "same values as in filter_ics r3014 (circa July 2007)" ;
data:

 MemberMetadata =
  "ensemble member      1",
  "ensemble member      2",
  "ensemble member      3",
  "ensemble member      4",
  "ensemble member      5",
  "ensemble member      6",
  "ensemble member      7",
  "ensemble member      8",
  "ensemble member      9",
  "ensemble member     10",
  "ensemble member     11",
  "ensemble member     12",
  "ensemble member     13",
  "ensemble member     14",
  "ensemble member     15",
  "ensemble member     16",
  "ensemble member     17",
  "ensemble member     18",
  "ensemble member     19",
  "ensemble member     20",
  "ensemble member     21",
  "ensemble member     22",
  "ensemble member     23",
  "ensemble member     24",
  "ensemble member     25",
  "ensemble member     26",
  "ensemble member     27",
  "ensemble member     28",
  "ensemble member     29",
  "ensemble member     30",
  "ensemble member     31",
  "ensemble member     32",
  "ensemble member     33",
  "ensemble member     34",
  "ensemble member     35",
  "ensemble member     36",
  "ensemble member     37",
  "ensemble member     38",
  "ensemble member     39",
  "ensemble member     40",
  "ensemble member     41",
  "ensemble member     42",
  "ensemble member     43",
  "ensemble member     44",
  "ensemble member     45",
  "ensemble member     46",
  "ensemble member     47",
  "ensemble member     48",
  "ensemble member     49",
  "ensemble member     50",
  "ensemble member     51",
  "ensemble member     52",
  "ensemble member     53",
  "ensemble member     54",
  "ensemble member     55",
  "ensemble member     56",
  "ensemble member     57",
  "ensemble member     58",
  "ensemble member     59",
  "ensemble member     60",
  "ensemble member     61",
  "ensemble member     62",
  "ensemble member     63",
  "ensemble member     64",
  "ensemble member     65",
  "ensemble member     66",
  "ensemble member     67",
  "ensemble member     68",
  "ensemble member     69",
  "ensemble member     70",
  "ensemble member     71",
  "ensemble member     72",
  "ensemble member     73",
  "ensemble member     74",
  "ensemble member     75",
  "ensemble member     76",
  "ensemble member     77",
  "ensemble member     78",
  "ensemble member     79",
  "ensemble member     80" ;

 concentration =
  5167.44927700767, 4479.15610033344, 5946.8985976654, 4880.76917157547, 
    7625.08271628216, 6154.93188217955, 5282.61877144751, 4471.73048833583, 
    3793.04031869691, 3094.91412937428,
  5071.41609860872, 4523.8939268231, 5963.43641555305, 4877.21878434774, 
    7589.91121070912, 6204.30508692013, 5367.3441052301, 4488.8592972656, 
    3745.80745869772, 3168.75038045218,
  5176.10965499913, 4526.62899442576, 5946.45733171349, 4912.63667707486, 
    7606.20912239408, 6181.68376525419, 5337.78620450484, 4456.98892091919, 
    3688.28100331018, 3126.76037132743,
  5147.14790191082, 4553.07313641949, 5951.9583612014, 4901.25848663976, 
    7586.94542964164, 6254.69698094819, 5366.26741644684, 4433.95779185845, 
    3817.52058398416, 3146.46889304371,
  5155.2952156588, 4471.53028354077, 5882.74349811162, 4992.93650256581, 
    7570.68953839956, 6172.59427395089, 5360.90746162091, 4455.52062380225, 
    3762.98202751411, 3129.78703203107,
  5081.81625347885, 4487.943124627, 5856.7237828836, 5005.12220790846, 
    7588.24938018252, 6204.15335330215, 5289.70532106749, 4427.44702762755, 
    3741.24984860258, 3165.44514826594,
  5147.88927786747, 4479.63167676891, 5915.36836685069, 4972.81610208727, 
    7555.07360459222, 6209.08910013202, 5309.92529979614, 4503.78393174698, 
    3735.40237088435, 3128.85111602778,
  5212.47544540583, 4522.72967728129, 5949.65153478115, 4906.69519268113, 
    7675.04081703867, 6142.21659859271, 5311.56873210376, 4471.55354626647, 
    3777.9901512883, 3094.67375377158,
  5201.55910863649, 4460.1750773373, 6061.40720499516, 4893.23401577366, 
    7655.7247612677, 6152.34038822817, 5360.81218728933, 4444.57387807784, 
    3773.76936773669, 3065.06651339611,
  5018.05951143294, 4501.58827460143, 5949.5208092236, 4883.14772223446, 
    7594.55345921469, 6168.20816590719, 5315.16580428916, 4466.99620335607, 
    3776.15182512405, 3105.20911679031,
  5139.87466886843, 4465.33660923562, 6006.44142737463, 4908.13733366068, 
    7590.15167600611, 6177.59653537969, 5363.99889406797, 4477.01957179019, 
    3751.03681235953, 3107.1644435788,
  5062.79553568938, 4551.84305292624, 5943.30565030342, 4913.66831743039, 
    7576.79605721191, 6186.55359421111, 5219.051439642, 4509.32807671859, 
    3769.38834988261, 3101.26300550372,
  5130.54216784188, 4480.44402009692, 5981.46783022331, 4892.51598116873, 
    7601.38688671873, 6192.21083215341, 5362.99845391557, 4497.62413671628, 
    3725.4059999813, 3167.74438128846,
  5190.71631245699, 4501.66611981571, 5999.50292491543, 4948.48060008286, 
    7533.76948597066, 6199.34795193482, 5350.92934593152, 4405.81306144864, 
    3792.89665623934, 3068.93386838865,
  5151.37116590051, 4542.31210721413, 5979.43422511503, 5015.08015252204, 
    7560.44275188729, 6221.21819130067, 5359.80950856632, 4387.7897403831, 
    3827.42821326138, 3145.70889778045,
  5155.25932821845, 4495.98684836379, 5965.89462808368, 4932.95687647224, 
    7516.87690217027, 6231.18368068678, 5293.48934158769, 4483.7767379716, 
    3754.68605652717, 3144.36189690583,
  5170.95715263564, 4494.28735699866, 5971.41999767849, 4940.68746151102, 
    7491.49760895883, 6216.57993064743, 5300.07081131948, 4499.76966064415, 
    3764.72212157166, 3124.31559784965,
  5074.71673877957, 4481.58387240951, 6008.23594718998, 4930.71510496826, 
    7708.83152093684, 6153.60583024395, 5294.9819577792, 4421.20248303127, 
    3771.65791288014, 3167.18285211219,
  5074.33074226474, 4538.62203343135, 5979.39702858008, 4932.94508484014, 
    7598.60093404636, 6224.92034715527, 5351.32025368635, 4445.90529105413, 
    3796.20717422531, 3106.50351920958,
  5063.81802297861, 4500.187175678, 5991.41005869297, 4987.25788033147, 
    7489.38505294453, 6166.22816661898, 5339.88477834268, 4438.64546829989, 
    3787.78587449296, 3131.64755875427,
  5167.80081323865, 4458.59003336545, 6025.13359522615, 4972.89494216159, 
    7575.72438067756, 6208.03993649735, 5282.11264349497, 4483.27871738451, 
    3675.72367172663, 3135.95217366964,
  5224.86605229394, 4494.02390424608, 6029.57654713715, 4993.27386319992, 
    7562.97465319504, 6212.98464885389, 5308.82353517207, 4491.79935463376, 
    3824.7615554802, 3115.12048563756,
  5099.96377460158, 4519.99702008152, 5924.07709229867, 4975.7632048603, 
    7555.02800031012, 6195.09300330218, 5341.33762199058, 4491.20357628811, 
    3768.70838777982, 3132.61559105481,
  5096.6543658565, 4502.06257594014, 6012.90884753178, 4898.99438294341, 
    7533.96989533136, 6261.15510774271, 5299.77309796176, 4412.6695412887, 
    3771.30948634677, 3118.15217726441,
  5137.15811290894, 4504.26369382418, 5969.59816441624, 5016.72596197525, 
    7511.10790774614, 6297.12394468955, 5269.98146193026, 4450.91964461768, 
    3719.81844835081, 3116.20152461885,
  5102.56580785841, 4549.11542804256, 5934.08105231417, 4932.20121554329, 
    7546.3587225934, 6177.32128288762, 5330.78952950057, 4441.54353754315, 
    3779.62466725837, 3192.41991368025,
  5150.99474723599, 4477.94798509355, 5947.5309284468, 4943.03212713642, 
    7601.53695495424, 6126.05727400066, 5292.18372531333, 4473.47835998095, 
    3791.48572565857, 3154.33161155157,
  5146.69877286376, 4480.50442308408, 5997.29223766494, 4936.66659107369, 
    7524.9053510833, 6189.0076085335, 5292.09356477614, 4493.63822392349, 
    3773.86606440472, 3175.15435199988,
  5141.90316997994, 4466.97945755218, 5973.46747599077, 4930.78837441487, 
    7533.33613505035, 6194.16128707273, 5355.64921338628, 4404.28314785369, 
    3780.59399738066, 3076.50272767856,
  5154.59139997614, 4445.58519116337, 5927.52433476045, 4939.18681305289, 
    7568.07923549269, 6235.45659919411, 5336.46302224864, 4518.29744224459, 
    3799.88700061455, 3102.42492108799,
  5070.64545145175, 4456.22249830144, 6033.11577308123, 4948.90435476985, 
    7625.2516449859, 6199.2902547825, 5323.77521449893, 4445.30140369698, 
    3779.23373869398, 3156.88239231121,
  5035.99368064126, 4516.0920733911, 5949.07685906715, 4949.39187967134, 
    7574.16490324597, 6268.72929766017, 5332.05787108937, 4422.89131413511, 
    3833.47622714989, 3169.1411539367,
  5151.9540963881, 4374.95072310076, 6049.18792682534, 4884.29192622718, 
    7618.69626356723, 6151.18102158092, 5376.43261798023, 4410.86796958741, 
    3754.1816589905, 3152.66039753779,
  5023.0261970124, 4464.98371503245, 5970.67175781262, 4968.24800583076, 
    7625.75915763929, 6223.40424865569, 5301.96150707024, 4450.73851484791, 
    3742.02986475977, 3121.83274726356,
  5113.64112532094, 4517.84097810781, 6007.70795284249, 4882.53223175353, 
    7661.39006469373, 6248.34723856012, 5279.02846521492, 4473.19756602326, 
    3735.74145851155, 3116.46620860281,
  5065.81073672435, 4515.53530920247, 5991.06374667026, 4919.61255696009, 
    7581.04486692895, 6260.28305365211, 5259.02964542701, 4475.32938552524, 
    3761.46688835003, 3178.16600581788,
  5083.24827026882, 4500.62017428399, 5859.48774972126, 5015.10551954802, 
    7442.57934776621, 6258.96895749554, 5312.66764332805, 4429.19305943997, 
    3775.20736740165, 3142.86231547555,
  5119.20023188893, 4512.16496945069, 5959.42864094804, 4926.64495901589, 
    7525.59843349722, 6222.12115941093, 5329.75286763736, 4452.39769427451, 
    3776.24548205451, 3162.25162112429,
  5164.87537740932, 4480.52155194355, 6004.09698917057, 4881.66020120269, 
    7669.27926172801, 6142.15575940293, 5366.90931309399, 4366.97177934759, 
    3840.58851120105, 3098.33685348768,
  5072.43575278185, 4508.01621246702, 5949.84961843017, 4925.21803553995, 
    7601.66879207006, 6177.54248527652, 5362.22328449341, 4436.53696829218, 
    3776.44347388997, 3151.20524122935,
  5083.78004523179, 4543.0135774296, 5963.53988292786, 4924.87556301359, 
    7543.98386703964, 6191.52023385607, 5333.7344274804, 4488.2494228577, 
    3727.77974395222, 3135.19431972596,
  5103.78358952497, 4513.70744846252, 5979.73844378255, 4990.51218893268, 
    7595.28784854708, 6196.55158240133, 5373.46541013225, 4456.06251847614, 
    3774.39492451967, 3097.15294523343,
  5086.62358697175, 4500.02750179481, 6002.2210661065, 4918.45414704982, 
    7585.11763998584, 6192.75337677432, 5369.36550635535, 4406.15418579766, 
    3757.91947788598, 3102.2194737499,
  5085.11173018242, 4428.78028087779, 6038.27480051974, 4889.66539165719, 
    7547.94675214865, 6161.39528160223, 5336.62077140202, 4435.54763263482, 
    3794.55484552035, 3123.03382634062,
  5150.02515183798, 4442.36410313491, 6022.57870123802, 4895.65042326048, 
    7619.27891721166, 6199.72648252036, 5324.601835837, 4453.4051265311, 
    3763.79472412435, 3182.93537278176,
  5140.74732963311, 4479.45856642697, 5918.72621144854, 4962.48528735283, 
    7523.63827920612, 6202.66707580731, 5344.80980364454, 4469.59270830628, 
    3834.76454088074, 3110.26862568632,
  5135.75599733995, 4516.98588660906, 5922.07852806346, 4906.26161793037, 
    7604.46740112674, 6115.92238312558, 5322.57979906159, 4447.53665341236, 
    3709.95947708309, 3143.0836650772,
  5148.50930807479, 4439.70642186281, 6035.50532204931, 4948.00373963122, 
    7491.55522343168, 6224.36247392485, 5299.52654200651, 4418.64979661556, 
    3724.79428725545, 3120.1369943302,
  5087.3217610848, 4453.89812134024, 6053.02411729208, 4894.01072171963, 
    7674.21464043177, 6155.85211470785, 5355.11888389967, 4478.61017509384, 
    3758.85576641768, 3129.02222966192,
  5101.03051062769, 4499.90122599631, 5918.05179036641, 4919.53336913724, 
    7664.87755108748, 6227.18734481841, 5264.59933557654, 4450.67895528259, 
    3808.60461554183, 3119.17645064334,
  5133.06995118887, 4480.77917842629, 6037.46953584176, 4928.52753863637, 
    7531.47756967442, 6188.01050823585, 5355.14577441995, 4436.54579339063, 
    3755.14677105684, 3157.48061356962,
  5115.28499388009, 4507.91717828197, 5945.13872201098, 4907.13971270896, 
    7668.71824343097, 6202.50818510863, 5309.81474867678, 4423.41789145573, 
    3738.5720258323, 3169.50745277754,
  5152.17427675414, 4518.76898521154, 6007.3017606535, 4924.86829426989, 
    7608.62532231945, 6183.07297045567, 5289.21966920952, 4498.49247407859, 
    3734.03398997481, 3193.16466907988,
  5194.70464102936, 4445.39617382015, 6014.94713580016, 4915.13583946702, 
    7569.46571799195, 6203.46238672913, 5230.83708825866, 4479.3261848975, 
    3820.25839907478, 3091.62167373297,
  5088.46226046481, 4523.00218889917, 5981.08730708784, 4895.33892337858, 
    7663.58359268814, 6180.8434363489, 5402.38853378578, 4440.35715835823, 
    3766.14983352117, 3181.14018132205,
  5153.35764870324, 4491.44927695577, 5994.73351970686, 4944.33002771072, 
    7622.16873317059, 6172.33931929537, 5368.63766107781, 4471.05842598785, 
    3729.24097415835, 3084.70112809135,
  5017.5647304342, 4465.19403102391, 6013.04128631556, 4957.23642705492, 
    7577.63129693762, 6167.4976184755, 5275.50242762597, 4462.74528873755, 
    3762.04185805478, 3156.22264886999,
  5106.86557068015, 4541.63579712852, 5935.13548564792, 4969.79469494356, 
    7559.03096175104, 6109.05682162077, 5355.12869963258, 4424.91993829343, 
    3760.28120607621, 3107.55808950264,
  5079.64096876566, 4540.16386421266, 6017.07435191535, 4858.80325960364, 
    7632.4762707954, 6210.14524229507, 5332.84645213476, 4449.20352088686, 
    3731.56600150898, 3110.21647828673,
  5101.95319503045, 4491.32585127161, 5996.70703261373, 4892.13931221763, 
    7647.09101920532, 6165.58531114141, 5343.83021641005, 4471.20916287605, 
    3720.95431471147, 3161.38643919079,
  5102.5273753359, 4494.27110082423, 5938.85824798176, 4894.62608052976, 
    7625.91741525265, 6166.58124268507, 5308.03832931209, 4419.48787558321, 
    3777.8197261267, 3155.58306928887,
  5173.76202474688, 4480.23358181992, 5956.1071021834, 4975.90484562343, 
    7628.74080700046, 6194.40268203292, 5348.25978604634, 4410.03915881923, 
    3791.91738760178, 3097.51716380827,
  5183.69807469949, 4463.55233060581, 5958.41163523256, 4975.34768621482, 
    7622.04379268469, 6206.41516390411, 5340.00730358964, 4492.71782343599, 
    3754.18535848988, 3052.85493041852,
  5132.81092778293, 4481.29333281875, 5943.49948355627, 4884.41117666636, 
    7641.92214408553, 6179.52175820595, 5316.20837605349, 4428.5421474545, 
    3744.82032132193, 3088.92132874764,
  5105.85949982479, 4510.66915670353, 5932.1521763856, 4969.44673466154, 
    7566.45701389151, 6200.92508630513, 5326.85297141165, 4400.01529165294, 
    3750.26512405343, 3181.24137933222,
  5148.05991180505, 4443.99193335487, 5956.4474458068, 4973.35084974135, 
    7585.11008200065, 6142.39655164642, 5345.96188209485, 4492.8683594801, 
    3693.16345784105, 3151.67759249838,
  5208.45107370593, 4490.32213043352, 5945.54777928061, 4963.3274564696, 
    7578.12753235643, 6188.87820725218, 5354.57277116957, 4443.05866961452, 
    3766.36361955924, 3099.88360386642,
  5115.84174527004, 4524.82199912879, 6043.9489622574, 4926.01283141416, 
    7504.73990426592, 6179.28068873198, 5351.21768259334, 4415.94801090923, 
    3766.00452067933, 3115.92619778007,
  5108.74567607368, 4502.63691228124, 6074.83191507215, 4940.10767003055, 
    7543.80202066171, 6204.77099906504, 5280.01429713246, 4460.01589209052, 
    3788.20368473418, 3165.72894027998,
  5032.33109445419, 4518.01455572718, 5933.3377263609, 4998.28942580928, 
    7517.23039099247, 6280.60146784494, 5351.37419154502, 4514.14234665451, 
    3775.42997470678, 3194.31368420811,
  5085.2153831422, 4491.54154747592, 5958.26624376263, 4901.65308259917, 
    7584.09417043027, 6176.42577525833, 5322.13161595452, 4513.30322913018, 
    3768.37107262586, 3140.11666197434,
  5103.59624065276, 4503.31334304895, 5869.26176369956, 4929.55013098015, 
    7484.19447738071, 6238.53641699289, 5315.29093956083, 4411.63497689205, 
    3765.10531492955, 3120.2718161626,
  5147.88589269751, 4480.47807173378, 5970.18423770196, 4925.35980334348, 
    7575.31514642887, 6206.27703742599, 5367.44456328351, 4462.27657317379, 
    3773.28319716578, 3132.23648282541,
  5063.7206543289, 4490.5112258112, 6036.41550057099, 4975.74101380984, 
    7507.85010458436, 6256.56801003897, 5297.74451449317, 4500.07536375217, 
    3728.5548182183, 3135.69638487578,
  5162.11774843347, 4457.20286528039, 6020.80214932017, 4893.06518672349, 
    7614.76390408391, 6164.15877305333, 5286.20692873376, 4469.78458188932, 
    3824.15261145156, 3042.04566991772,
  5039.39010303376, 4506.79447991978, 6004.03728040389, 4946.22877244145, 
    7604.26979889153, 6151.04558111486, 5349.2625075676, 4492.05937721383, 
    3777.77360522594, 3119.78489566798,
  5191.94892030821, 4482.70603287449, 5952.15603201574, 4953.51971071743, 
    7513.2929722302, 6308.41666987499, 5272.32177279519, 4443.17624568108, 
    3748.21415231144, 3096.18228868378,
  5093.89203400228, 4512.67304659479, 5928.46862995695, 4919.06050721316, 
    7508.15594832963, 6274.83022561345, 5357.42153730051, 4463.81143583754, 
    3809.13354055303, 3112.81843383716,
  5118.39724821137, 4494.56820491257, 5988.19905472261, 4998.83631972666, 
    7564.55337256294, 6240.38520293211, 5304.35181352085, 4526.53579316383, 
    3782.81207673978, 3131.3581184442,
  5068.66047927635, 4493.81790520062, 5957.69205397143, 4946.15856801485, 
    7596.22433577696, 6097.3978846894, 5383.98998392653, 4447.76157704973, 
    3739.15692835372, 3151.08492992999 ;

 mean_source =
  0.9999999999999, 0.0999999999999897, 0.9999999999999, 0.0999999999999897, 
    0.9999999999999, 0.0999999999999897, 0.0999999999999897, 
    0.0999999999999897, 0.0999999999999897, 0.0999999999999897,
  0.999999999999804, 0.0999999999999801, 0.999999999999804, 
    0.0999999999999801, 0.999999999999804, 0.0999999999999801, 
    0.0999999999999801, 0.0999999999999801, 0.0999999999999801, 
    0.0999999999999801,
  0.999999999999947, 0.0999999999999945, 0.999999999999947, 
    0.0999999999999945, 0.999999999999947, 0.0999999999999945, 
    0.0999999999999945, 0.0999999999999945, 0.0999999999999945, 
    0.0999999999999945,
  0.999999999999755, 0.0999999999999752, 0.999999999999755, 
    0.0999999999999752, 0.999999999999755, 0.0999999999999752, 
    0.0999999999999752, 0.0999999999999752, 0.0999999999999752, 
    0.0999999999999752,
  0.999999999999978, 0.0999999999999975, 0.999999999999978, 
    0.0999999999999975, 0.999999999999978, 0.0999999999999975, 
    0.0999999999999975, 0.0999999999999975, 0.0999999999999975, 
    0.0999999999999975,
  1.0000000000001, 0.10000000000001, 1.0000000000001, 0.10000000000001, 
    1.0000000000001, 0.10000000000001, 0.10000000000001, 0.10000000000001, 
    0.10000000000001, 0.10000000000001,
  1.00000000000006, 0.100000000000005, 1.00000000000006, 0.100000000000005, 
    1.00000000000006, 0.100000000000005, 0.100000000000005, 
    0.100000000000005, 0.100000000000005, 0.100000000000005,
  0.999999999999816, 0.0999999999999813, 0.999999999999816, 
    0.0999999999999813, 0.999999999999816, 0.0999999999999813, 
    0.0999999999999813, 0.0999999999999813, 0.0999999999999813, 
    0.0999999999999813,
  0.999999999999858, 0.0999999999999854, 0.999999999999858, 
    0.0999999999999854, 0.999999999999858, 0.0999999999999854, 
    0.0999999999999854, 0.0999999999999854, 0.0999999999999854, 
    0.0999999999999854,
  0.999999999999799, 0.0999999999999797, 0.999999999999799, 
    0.0999999999999797, 0.999999999999799, 0.0999999999999797, 
    0.0999999999999797, 0.0999999999999797, 0.0999999999999797, 
    0.0999999999999797,
  0.99999999999973, 0.0999999999999728, 0.99999999999973, 0.0999999999999728, 
    0.99999999999973, 0.0999999999999728, 0.0999999999999728, 
    0.0999999999999728, 0.0999999999999728, 0.0999999999999728,
  0.99999999999991, 0.0999999999999907, 0.99999999999991, 0.0999999999999907, 
    0.99999999999991, 0.0999999999999907, 0.0999999999999907, 
    0.0999999999999907, 0.0999999999999907, 0.0999999999999907,
  0.999999999999868, 0.0999999999999864, 0.999999999999868, 
    0.0999999999999864, 0.999999999999868, 0.0999999999999864, 
    0.0999999999999864, 0.0999999999999864, 0.0999999999999864, 
    0.0999999999999864,
  0.99999999999991, 0.0999999999999907, 0.99999999999991, 0.0999999999999907, 
    0.99999999999991, 0.0999999999999907, 0.0999999999999907, 
    0.0999999999999907, 0.0999999999999907, 0.0999999999999907,
  0.999999999999874, 0.099999999999987, 0.999999999999874, 0.099999999999987, 
    0.999999999999874, 0.099999999999987, 0.099999999999987, 
    0.099999999999987, 0.099999999999987, 0.099999999999987,
  1.00000000000001, 0.1, 1.00000000000001, 0.1, 1.00000000000001, 0.1, 0.1, 
    0.1, 0.1, 0.1,
  0.999999999999749, 0.0999999999999746, 0.999999999999749, 
    0.0999999999999746, 0.999999999999749, 0.0999999999999746, 
    0.0999999999999746, 0.0999999999999746, 0.0999999999999746, 
    0.0999999999999746,
  0.999999999999946, 0.0999999999999941, 0.999999999999946, 
    0.0999999999999941, 0.999999999999946, 0.0999999999999941, 
    0.0999999999999941, 0.0999999999999941, 0.0999999999999941, 
    0.0999999999999941,
  0.999999999999838, 0.0999999999999836, 0.999999999999838, 
    0.0999999999999836, 0.999999999999838, 0.0999999999999836, 
    0.0999999999999836, 0.0999999999999836, 0.0999999999999836, 
    0.0999999999999836,
  0.999999999999747, 0.0999999999999744, 0.999999999999747, 
    0.0999999999999744, 0.999999999999747, 0.0999999999999744, 
    0.0999999999999744, 0.0999999999999744, 0.0999999999999744, 
    0.0999999999999744,
  0.999999999999856, 0.0999999999999853, 0.999999999999856, 
    0.0999999999999853, 0.999999999999856, 0.0999999999999853, 
    0.0999999999999853, 0.0999999999999853, 0.0999999999999853, 
    0.0999999999999853,
  0.999999999999899, 0.0999999999999895, 0.999999999999899, 
    0.0999999999999895, 0.999999999999899, 0.0999999999999895, 
    0.0999999999999895, 0.0999999999999895, 0.0999999999999895, 
    0.0999999999999895,
  0.99999999999981, 0.0999999999999807, 0.99999999999981, 0.0999999999999807, 
    0.99999999999981, 0.0999999999999807, 0.0999999999999807, 
    0.0999999999999807, 0.0999999999999807, 0.0999999999999807,
  0.999999999999771, 0.0999999999999767, 0.999999999999771, 
    0.0999999999999767, 0.999999999999771, 0.0999999999999767, 
    0.0999999999999767, 0.0999999999999767, 0.0999999999999767, 
    0.0999999999999767,
  0.99999999999994, 0.0999999999999936, 0.99999999999994, 0.0999999999999936, 
    0.99999999999994, 0.0999999999999936, 0.0999999999999936, 
    0.0999999999999936, 0.0999999999999936, 0.0999999999999936,
  0.999999999999975, 0.0999999999999973, 0.999999999999975, 
    0.0999999999999973, 0.999999999999975, 0.0999999999999973, 
    0.0999999999999973, 0.0999999999999973, 0.0999999999999973, 
    0.0999999999999973,
  0.999999999999838, 0.0999999999999835, 0.999999999999838, 
    0.0999999999999835, 0.999999999999838, 0.0999999999999835, 
    0.0999999999999835, 0.0999999999999835, 0.0999999999999835, 
    0.0999999999999835,
  0.999999999999774, 0.0999999999999771, 0.999999999999774, 
    0.0999999999999771, 0.999999999999774, 0.0999999999999771, 
    0.0999999999999771, 0.0999999999999771, 0.0999999999999771, 
    0.0999999999999771,
  0.999999999999811, 0.099999999999981, 0.999999999999811, 0.099999999999981, 
    0.999999999999811, 0.099999999999981, 0.099999999999981, 
    0.099999999999981, 0.099999999999981, 0.099999999999981,
  0.999999999999969, 0.0999999999999965, 0.999999999999969, 
    0.0999999999999965, 0.999999999999969, 0.0999999999999965, 
    0.0999999999999965, 0.0999999999999965, 0.0999999999999965, 
    0.0999999999999965,
  0.999999999999941, 0.0999999999999938, 0.999999999999941, 
    0.0999999999999938, 0.999999999999941, 0.0999999999999938, 
    0.0999999999999938, 0.0999999999999938, 0.0999999999999938, 
    0.0999999999999938,
  1.00000000000002, 0.100000000000002, 1.00000000000002, 0.100000000000002, 
    1.00000000000002, 0.100000000000002, 0.100000000000002, 
    0.100000000000002, 0.100000000000002, 0.100000000000002,
  1.00000000000011, 0.10000000000001, 1.00000000000011, 0.10000000000001, 
    1.00000000000011, 0.10000000000001, 0.10000000000001, 0.10000000000001, 
    0.10000000000001, 0.10000000000001,
  0.999999999999738, 0.0999999999999735, 0.999999999999738, 
    0.0999999999999735, 0.999999999999738, 0.0999999999999735, 
    0.0999999999999735, 0.0999999999999735, 0.0999999999999735, 
    0.0999999999999735,
  1.00000000000006, 0.100000000000005, 1.00000000000006, 0.100000000000005, 
    1.00000000000006, 0.100000000000005, 0.100000000000005, 
    0.100000000000005, 0.100000000000005, 0.100000000000005,
  1.00000000000002, 0.100000000000002, 1.00000000000002, 0.100000000000002, 
    1.00000000000002, 0.100000000000002, 0.100000000000002, 
    0.100000000000002, 0.100000000000002, 0.100000000000002,
  0.999999999999922, 0.0999999999999919, 0.999999999999922, 
    0.0999999999999919, 0.999999999999922, 0.0999999999999919, 
    0.0999999999999919, 0.0999999999999919, 0.0999999999999919, 
    0.0999999999999919,
  0.999999999999838, 0.0999999999999835, 0.999999999999838, 
    0.0999999999999835, 0.999999999999838, 0.0999999999999835, 
    0.0999999999999835, 0.0999999999999835, 0.0999999999999835, 
    0.0999999999999835,
  0.999999999999926, 0.0999999999999922, 0.999999999999926, 
    0.0999999999999922, 0.999999999999926, 0.0999999999999922, 
    0.0999999999999922, 0.0999999999999922, 0.0999999999999922, 
    0.0999999999999922,
  1.00000000000004, 0.100000000000004, 1.00000000000004, 0.100000000000004, 
    1.00000000000004, 0.100000000000004, 0.100000000000004, 
    0.100000000000004, 0.100000000000004, 0.100000000000004,
  1.00000000000013, 0.100000000000013, 1.00000000000013, 0.100000000000013, 
    1.00000000000013, 0.100000000000013, 0.100000000000013, 
    0.100000000000013, 0.100000000000013, 0.100000000000013,
  0.999999999999893, 0.0999999999999889, 0.999999999999893, 
    0.0999999999999889, 0.999999999999893, 0.0999999999999889, 
    0.0999999999999889, 0.0999999999999889, 0.0999999999999889, 
    0.0999999999999889,
  0.999999999999942, 0.0999999999999941, 0.999999999999942, 
    0.0999999999999941, 0.999999999999942, 0.0999999999999941, 
    0.0999999999999941, 0.0999999999999941, 0.0999999999999941, 
    0.0999999999999941,
  0.999999999999725, 0.0999999999999722, 0.999999999999725, 
    0.0999999999999722, 0.999999999999725, 0.0999999999999722, 
    0.0999999999999722, 0.0999999999999722, 0.0999999999999722, 
    0.0999999999999722,
  0.999999999999721, 0.0999999999999719, 0.999999999999721, 
    0.0999999999999719, 0.999999999999721, 0.0999999999999719, 
    0.0999999999999719, 0.0999999999999719, 0.0999999999999719, 
    0.0999999999999719,
  0.999999999999729, 0.0999999999999725, 0.999999999999729, 
    0.0999999999999725, 0.999999999999729, 0.0999999999999725, 
    0.0999999999999725, 0.0999999999999725, 0.0999999999999725, 
    0.0999999999999725,
  0.999999999999847, 0.0999999999999843, 0.999999999999847, 
    0.0999999999999843, 0.999999999999847, 0.0999999999999843, 
    0.0999999999999843, 0.0999999999999843, 0.0999999999999843, 
    0.0999999999999843,
  0.999999999999907, 0.0999999999999904, 0.999999999999907, 
    0.0999999999999904, 0.999999999999907, 0.0999999999999904, 
    0.0999999999999904, 0.0999999999999904, 0.0999999999999904, 
    0.0999999999999904,
  0.999999999999812, 0.0999999999999808, 0.999999999999812, 
    0.0999999999999808, 0.999999999999812, 0.0999999999999808, 
    0.0999999999999808, 0.0999999999999808, 0.0999999999999808, 
    0.0999999999999808,
  0.99999999999966, 0.0999999999999657, 0.99999999999966, 0.0999999999999657, 
    0.99999999999966, 0.0999999999999657, 0.0999999999999657, 
    0.0999999999999657, 0.0999999999999657, 0.0999999999999657,
  0.999999999999782, 0.0999999999999778, 0.999999999999782, 
    0.0999999999999778, 0.999999999999782, 0.0999999999999778, 
    0.0999999999999778, 0.0999999999999778, 0.0999999999999778, 
    0.0999999999999778,
  0.999999999999943, 0.0999999999999942, 0.999999999999943, 
    0.0999999999999942, 0.999999999999943, 0.0999999999999942, 
    0.0999999999999942, 0.0999999999999942, 0.0999999999999942, 
    0.0999999999999942,
  0.999999999999883, 0.099999999999988, 0.999999999999883, 0.099999999999988, 
    0.999999999999883, 0.099999999999988, 0.099999999999988, 
    0.099999999999988, 0.099999999999988, 0.099999999999988,
  0.999999999999965, 0.0999999999999962, 0.999999999999965, 
    0.0999999999999962, 0.999999999999965, 0.0999999999999962, 
    0.0999999999999962, 0.0999999999999962, 0.0999999999999962, 
    0.0999999999999962,
  0.999999999999922, 0.0999999999999917, 0.999999999999922, 
    0.0999999999999917, 0.999999999999922, 0.0999999999999917, 
    0.0999999999999917, 0.0999999999999917, 0.0999999999999917, 
    0.0999999999999917,
  0.999999999999911, 0.0999999999999908, 0.999999999999911, 
    0.0999999999999908, 0.999999999999911, 0.0999999999999908, 
    0.0999999999999908, 0.0999999999999908, 0.0999999999999908, 
    0.0999999999999908,
  0.999999999999845, 0.0999999999999841, 0.999999999999845, 
    0.0999999999999841, 0.999999999999845, 0.0999999999999841, 
    0.0999999999999841, 0.0999999999999841, 0.0999999999999841, 
    0.0999999999999841,
  0.999999999999656, 0.0999999999999652, 0.999999999999656, 
    0.0999999999999652, 0.999999999999656, 0.0999999999999652, 
    0.0999999999999652, 0.0999999999999652, 0.0999999999999652, 
    0.0999999999999652,
  0.999999999999809, 0.0999999999999806, 0.999999999999809, 
    0.0999999999999806, 0.999999999999809, 0.0999999999999806, 
    0.0999999999999806, 0.0999999999999806, 0.0999999999999806, 
    0.0999999999999806,
  1.00000000000005, 0.100000000000005, 1.00000000000005, 0.100000000000005, 
    1.00000000000005, 0.100000000000005, 0.100000000000005, 
    0.100000000000005, 0.100000000000005, 0.100000000000005,
  0.999999999999919, 0.0999999999999916, 0.999999999999919, 
    0.0999999999999916, 0.999999999999919, 0.0999999999999916, 
    0.0999999999999916, 0.0999999999999916, 0.0999999999999916, 
    0.0999999999999916,
  0.999999999999944, 0.0999999999999941, 0.999999999999944, 
    0.0999999999999941, 0.999999999999944, 0.0999999999999941, 
    0.0999999999999941, 0.0999999999999941, 0.0999999999999941, 
    0.0999999999999941,
  0.99999999999992, 0.0999999999999916, 0.99999999999992, 0.0999999999999916, 
    0.99999999999992, 0.0999999999999916, 0.0999999999999916, 
    0.0999999999999916, 0.0999999999999916, 0.0999999999999916,
  1.00000000000013, 0.100000000000012, 1.00000000000013, 0.100000000000012, 
    1.00000000000013, 0.100000000000012, 0.100000000000012, 
    0.100000000000012, 0.100000000000012, 0.100000000000012,
  0.999999999999861, 0.0999999999999858, 0.999999999999861, 
    0.0999999999999858, 0.999999999999861, 0.0999999999999858, 
    0.0999999999999858, 0.0999999999999858, 0.0999999999999858, 
    0.0999999999999858,
  0.999999999999713, 0.099999999999971, 0.999999999999713, 0.099999999999971, 
    0.999999999999713, 0.099999999999971, 0.099999999999971, 
    0.099999999999971, 0.099999999999971, 0.099999999999971,
  0.999999999999789, 0.0999999999999786, 0.999999999999789, 
    0.0999999999999786, 0.999999999999789, 0.0999999999999786, 
    0.0999999999999786, 0.0999999999999786, 0.0999999999999786, 
    0.0999999999999786,
  1.00000000000002, 0.100000000000002, 1.00000000000002, 0.100000000000002, 
    1.00000000000002, 0.100000000000002, 0.100000000000002, 
    0.100000000000002, 0.100000000000002, 0.100000000000002,
  0.999999999999827, 0.0999999999999824, 0.999999999999827, 
    0.0999999999999824, 0.999999999999827, 0.0999999999999824, 
    0.0999999999999824, 0.0999999999999824, 0.0999999999999824, 
    0.0999999999999824,
  0.999999999999766, 0.0999999999999763, 0.999999999999766, 
    0.0999999999999763, 0.999999999999766, 0.0999999999999763, 
    0.0999999999999763, 0.0999999999999763, 0.0999999999999763, 
    0.0999999999999763,
  0.999999999999708, 0.0999999999999705, 0.999999999999708, 
    0.0999999999999705, 0.999999999999708, 0.0999999999999705, 
    0.0999999999999705, 0.0999999999999705, 0.0999999999999705, 
    0.0999999999999705,
  0.99999999999981, 0.0999999999999805, 0.99999999999981, 0.0999999999999805, 
    0.99999999999981, 0.0999999999999805, 0.0999999999999805, 
    0.0999999999999805, 0.0999999999999805, 0.0999999999999805,
  0.999999999999792, 0.0999999999999788, 0.999999999999792, 
    0.0999999999999788, 0.999999999999792, 0.0999999999999788, 
    0.0999999999999788, 0.0999999999999788, 0.0999999999999788, 
    0.0999999999999788,
  0.999999999999968, 0.0999999999999965, 0.999999999999968, 
    0.0999999999999965, 0.999999999999968, 0.0999999999999965, 
    0.0999999999999965, 0.0999999999999965, 0.0999999999999965, 
    0.0999999999999965,
  0.999999999999808, 0.0999999999999804, 0.999999999999808, 
    0.0999999999999804, 0.999999999999808, 0.0999999999999804, 
    0.0999999999999804, 0.0999999999999804, 0.0999999999999804, 
    0.0999999999999804,
  1.00000000000009, 0.100000000000009, 1.00000000000009, 0.100000000000009, 
    1.00000000000009, 0.100000000000009, 0.100000000000009, 
    0.100000000000009, 0.100000000000009, 0.100000000000009,
  0.999999999999861, 0.0999999999999858, 0.999999999999861, 
    0.0999999999999858, 0.999999999999861, 0.0999999999999858, 
    0.0999999999999858, 0.0999999999999858, 0.0999999999999858, 
    0.0999999999999858,
  0.999999999999852, 0.0999999999999848, 0.999999999999852, 
    0.0999999999999848, 0.999999999999852, 0.0999999999999848, 
    0.0999999999999848, 0.0999999999999848, 0.0999999999999848, 
    0.0999999999999848,
  1.00000000000001, 0.100000000000001, 1.00000000000001, 0.100000000000001, 
    1.00000000000001, 0.100000000000001, 0.100000000000001, 
    0.100000000000001, 0.100000000000001, 0.100000000000001,
  0.999999999999839, 0.0999999999999835, 0.999999999999839, 
    0.0999999999999835, 0.999999999999839, 0.0999999999999835, 
    0.0999999999999835, 0.0999999999999835, 0.0999999999999835, 
    0.0999999999999835 ;

 source =
  0.705066638243117, 0.0733340783104723, 0.629917887536483, 
    0.0332779173368713, 1.04919926460651, 0.0770801224980458, 
    0.11212832381492, 0.0546879329523612, 0.0891561839104128, 
    0.0795008330231803,
  0.589834972600891, 0.107892707559408, 0.596778933105225, 
    0.0419081069304474, 1.12344811523075, 0.0681109153960028, 
    0.138533647187574, 0.0758994021291895, 0.0928349547795532, 
    0.096602369335389,
  0.681827846284297, 0.0967325331958445, 0.600887945000227, 
    0.0569527603893311, 0.974154309825333, 0.0672536388164413, 
    0.124525603112663, 0.0798412590077007, 0.0732096948567109, 
    0.100535888860457,
  0.765745788553062, 0.102382827048167, 0.648388167236289, 
    0.0559688842675797, 1.18249454566717, 0.0703225538836658, 
    0.112694065311461, 0.0654023766261767, 0.0864067149859118, 
    0.0902174196800763,
  0.676400875097642, 0.106410931075695, 0.643349740871845, 
    0.0655635512665382, 1.08129435252258, 0.0897419253004563, 
    0.131239123951426, 0.0753161139307684, 0.07833780617769, 
    0.0831192225731204,
  0.622378774563618, 0.11695928685218, 0.579940717154545, 0.060498837406311, 
    1.0588182911002, 0.0810792926441456, 0.122713086262476, 
    0.0689879503920323, 0.0791092753776901, 0.0916632962128114,
  0.671956773198338, 0.0910038366567827, 0.63343896886984, 
    0.0477398878090905, 1.05640465212531, 0.0673989707832787, 
    0.121965664953757, 0.0752153192683271, 0.0796158610161598, 
    0.103130406919556,
  0.620712314922599, 0.112473131382374, 0.638700306482544, 
    0.0397894653611385, 1.06714106398264, 0.0685622013987092, 
    0.120777671644203, 0.0639207706331109, 0.0970714648437485, 
    0.0838870007424036,
  0.689438762727159, 0.0927472424325867, 0.695120117324176, 
    0.0442582270987189, 1.07699197630329, 0.0758101876381765, 
    0.132428659318116, 0.0472598832144668, 0.0826855988361657, 
    0.096616054386262,
  0.680049176045974, 0.110461270970457, 0.607617367181005, 
    0.0443740234162227, 1.03374566773973, 0.0689303293807305, 
    0.133263135707944, 0.0603578890389959, 0.0972937051743012, 
    0.0736913242289614,
  0.711042976470512, 0.0907659444101589, 0.676193668198507, 
    0.0511987209679455, 0.994126443761716, 0.0843522170825941, 
    0.11585909989878, 0.0648306779179122, 0.0676712729061231, 
    0.0889977554596593,
  0.610146998181197, 0.100511249510745, 0.599713373870491, 
    0.0502465414054797, 1.13716094408766, 0.0703087698840655, 
    0.124798635973711, 0.0619727660837626, 0.0844072318170184, 
    0.0824562549540519,
  0.674250099957889, 0.107516989614221, 0.64554388401195, 0.0675983824763516, 
    1.12159933757059, 0.0801532284789292, 0.11861758537113, 
    0.0688749232006998, 0.0739362991406229, 0.101417137131104,
  0.760731379814478, 0.11634379296338, 0.638042587089311, 0.0551056484531637, 
    1.02259688170265, 0.0773568853017502, 0.137755336538072, 
    0.0830541243956231, 0.0786677135505595, 0.0795800453291728,
  0.640962184671513, 0.0957953912155348, 0.617259348825695, 
    0.0537312165033953, 0.973592740059966, 0.0695755727375122, 
    0.133746712390475, 0.0587486702407893, 0.0935420497163756, 
    0.087676676964408,
  0.66082862419894, 0.0852422489521663, 0.640811369595745, 
    0.0488880967474506, 0.989408397703155, 0.0811855121436139, 
    0.122024886976145, 0.0665418972668005, 0.0997287764566224, 
    0.0988334027426457,
  0.643113126548904, 0.100748230442888, 0.644607003645239, 
    0.0672987280302069, 1.09280405599085, 0.0698301238646935, 
    0.108302210378581, 0.0705140904392185, 0.0837851146840673, 
    0.0777627806449251,
  0.682704468869028, 0.0833857396500958, 0.641250595267399, 
    0.0320341198664644, 1.07159876650734, 0.0501559380740376, 
    0.120059024511505, 0.0550079044258249, 0.0980049310352754, 
    0.0982007533253182,
  0.617864279589507, 0.0938290965701267, 0.63215982336708, 
    0.0556858241663058, 1.04360781394016, 0.0498357939098701, 
    0.133814507796847, 0.060699394625236, 0.0979785581590735, 
    0.0803011871300926,
  0.662659399276336, 0.106458750152749, 0.700511952191131, 
    0.0425319168039038, 1.01298274779164, 0.0717090112391603, 
    0.126979150309721, 0.0599590691446759, 0.0816128584568972, 
    0.0917086285012759,
  0.645654018171173, 0.0965701729821541, 0.634700945821621, 
    0.0458237099369291, 1.06946433122064, 0.0759142349148394, 
    0.109287896873288, 0.052484410508573, 0.0680059028785863, 
    0.092898828602115,
  0.7082647062345, 0.0979565220065729, 0.684815846749953, 0.0474609935341565, 
    1.040175439079, 0.0802406733551489, 0.126455402357598, 
    0.0682947113911633, 0.0955756794258996, 0.0852725688786577,
  0.662950887561494, 0.0905160886384081, 0.691912596774246, 
    0.0468461840526323, 1.08657085708293, 0.0655101928925995, 
    0.133181099897822, 0.0609114761224656, 0.0837776903219462, 
    0.0916615454628122,
  0.620384429174498, 0.108892552101973, 0.660602345197835, 
    0.0453086292345544, 1.0654127421779, 0.0767709640764224, 
    0.129819297031361, 0.0644056473974526, 0.0764119380717949, 
    0.0876315473662141,
  0.689758757764923, 0.0979866010962744, 0.642002235614288, 
    0.0437484729488665, 1.01616730297991, 0.0837304478408763, 
    0.119529921359897, 0.0635826020027, 0.0782364148478441, 0.0759685312774835,
  0.635673054508252, 0.0985021687599732, 0.625610821149025, 
    0.044739687054915, 1.05297641704805, 0.0768216054505485, 
    0.133382466399506, 0.0712045289266711, 0.0977988357232542, 
    0.0980731154183136,
  0.669751906206873, 0.112205326849118, 0.621822780530661, 
    0.0513881943664011, 0.980926902566055, 0.0775016374423663, 
    0.13183218895439, 0.0716146258874958, 0.0918339362011841, 
    0.0915085206427916,
  0.712053956319683, 0.0977298910252042, 0.567238734120884, 
    0.0482848022653349, 1.08612228933093, 0.0657681404733733, 
    0.111682239441401, 0.0747568549526846, 0.0688725470124708, 
    0.092708181310192,
  0.659359621683122, 0.0956694836154842, 0.632884943120326, 
    0.0532154840201283, 1.12185126022191, 0.0642003920221279, 
    0.132984808550129, 0.0577551884230839, 0.102677213251034, 
    0.0994912539363729,
  0.687979670310914, 0.0891821375924655, 0.593460355154029, 
    0.0289027995636321, 1.11438931772824, 0.077734813045509, 
    0.126637301685775, 0.0669597209758471, 0.0849433896576314, 
    0.0833742618586422,
  0.698825646419242, 0.0902347129372859, 0.678144923074957, 
    0.0539060203095569, 1.05560590821445, 0.0724236031069346, 
    0.133475887591415, 0.0496684284360892, 0.0776260648391858, 
    0.0986589516061716,
  0.5950712038126, 0.103196722863574, 0.58417087530365, 0.0584002723141047, 
    1.04748499274646, 0.0580370186848278, 0.132465909002187, 
    0.0520887297494337, 0.0925808744008971, 0.0917295347090934,
  0.6011242847305, 0.0949575390245851, 0.692069562915291, 0.0646437015679463, 
    0.971936382782245, 0.0779328143766433, 0.137435662966023, 
    0.0509785954418866, 0.0858880167987677, 0.0947239210984222,
  0.601311665023304, 0.101977268558375, 0.605099042798309, 
    0.0394971601260537, 1.06868693517197, 0.0797861980359071, 
    0.123244473483407, 0.0876836646287271, 0.0889134055440988, 
    0.0929666422876467,
  0.648608371993195, 0.109087768791199, 0.58820918664395, 0.055695844266555, 
    1.1202609184884, 0.0781314825276315, 0.124733392804091, 
    0.0646486311275935, 0.0841443381463957, 0.0988732274035227,
  0.722159151727599, 0.123801297171799, 0.671626574261902, 
    0.0662405771387729, 1.05758201501465, 0.0905156152746159, 
    0.116962344016812, 0.087326137819114, 0.0818051160095755, 
    0.109172536479204,
  0.66409856232126, 0.097292720799141, 0.632000874428786, 0.0488816377293866, 
    1.03788580786798, 0.0792945173620004, 0.117036524455902, 
    0.0563187997211358, 0.0920085127279908, 0.103995960244487,
  0.678236634393544, 0.107497041565445, 0.66792268004384, 0.0697633859737304, 
    1.01858824719267, 0.0791683829780354, 0.112438211629884, 
    0.0669294174974982, 0.097966234028533, 0.0954182091909361,
  0.626142122488711, 0.107138401203267, 0.636015707902463, 
    0.0444954046697436, 1.1017180132622, 0.0647439377689195, 
    0.134769386577317, 0.0553639405399374, 0.105436015216114, 
    0.085441202731971,
  0.671891102525808, 0.115227919545619, 0.608958256182995, 
    0.0428784462795609, 1.13867010525082, 0.0660880798312595, 
    0.126800358027802, 0.061580330527744, 0.0815512206011445, 
    0.100614151599338,
  0.650282950140716, 0.098014399145221, 0.662119008963061, 
    0.0501130555106218, 1.0166757368047, 0.0677982949986168, 
    0.127164870976532, 0.0500087949592818, 0.0919013597546026, 
    0.105555419061003,
  0.678238690235669, 0.101127146546573, 0.637511976916254, 
    0.0591302553461783, 1.07076989970187, 0.0856172349071454, 
    0.114043731093709, 0.0847399371279573, 0.100941840365796, 
    0.0786605615920374,
  0.663345062726248, 0.0950219584993322, 0.691457952559562, 
    0.0643080141041463, 1.13416147859567, 0.0708016876650868, 
    0.139086399322518, 0.0695336602974748, 0.0872703256835945, 
    0.0865598927256709,
  0.652154557258634, 0.0925862762712977, 0.630655294176615, 
    0.0514171990564296, 1.06710518776796, 0.0781263385052347, 
    0.120106415083641, 0.0695971563616093, 0.104784215258485, 
    0.0825523997972238,
  0.606473033845002, 0.0912019384899658, 0.692805826713699, 
    0.0408187163130568, 1.01353519941901, 0.0814336167284537, 
    0.12725888418972, 0.0682536321903201, 0.094406966780556, 
    0.0897400759425526,
  0.687911062266219, 0.100024027112243, 0.658122896752907, 
    0.0528449112506048, 1.02084871465884, 0.0537337738145384, 
    0.139033992132066, 0.0537541591925158, 0.103104954004018, 
    0.0714231284978951,
  0.690073754238752, 0.110736855045154, 0.607255111040356, 
    0.0578866582023021, 0.981785584223066, 0.0758200994167771, 
    0.124162997208306, 0.0670231061052974, 0.0752750509089051, 
    0.0904421059920949,
  0.688959430213984, 0.0727036220630946, 0.632157581735596, 
    0.0414302194105534, 1.14414144110721, 0.0742763134169771, 
    0.117294804810063, 0.0547417768089816, 0.0887766275192507, 
    0.0818435013942807,
  0.570495242526084, 0.102266179730857, 0.646303969622987, 
    0.0514253434405374, 1.08900792875935, 0.0751088634856464, 
    0.12047123446746, 0.0513390997370826, 0.0857986398165543, 
    0.0863803357104582,
  0.664777039206035, 0.0934939715456683, 0.612046256279605, 
    0.0599326029387711, 1.06207567360342, 0.0802350492750331, 
    0.124070297136299, 0.0666635497183775, 0.0854480548137757, 
    0.0938044763297795,
  0.654077693907151, 0.117362602680891, 0.553277178030285, 
    0.0472299820687585, 1.09915783818572, 0.0698234937548714, 
    0.141080646724261, 0.0740753174100979, 0.083026948925883, 
    0.0919443417226003,
  0.68910451512705, 0.100822922398259, 0.658704909634032, 0.0476402338898636, 
    1.024820985024, 0.0609319279270842, 0.1143450000624, 0.0605942365060833, 
    0.073236528403639, 0.0944354557441919,
  0.70345776674289, 0.0933971733755828, 0.640323613998067, 
    0.0662316729833076, 1.07841287856021, 0.0840766141675628, 
    0.118787265134419, 0.0687893606912623, 0.0738050263672607, 
    0.0944398940981504,
  0.68859714984435, 0.0807031857828808, 0.570082665977144, 
    0.0429438167495444, 1.07578843373538, 0.06953671482474, 
    0.112698883597915, 0.0766784778530921, 0.0861983676179856, 
    0.0830384802556754,
  0.740671668770105, 0.0923529124867053, 0.634287354982064, 
    0.0489651872525976, 1.09037250877955, 0.0796240192391989, 
    0.119998038543379, 0.0515435168492264, 0.0740379486577101, 
    0.086032746737788,
  0.656189723930539, 0.111823066083333, 0.617165983187478, 0.046707917015552, 
    1.02603742595306, 0.0777275170324892, 0.141360657121012, 
    0.0790263843621564, 0.0829771604642023, 0.1031916310453,
  0.637264126763233, 0.0939091298411044, 0.6333032053021, 0.0712750950853702, 
    1.00429759695573, 0.0815096567516702, 0.115171453578749, 
    0.0731155443305133, 0.068649968363095, 0.0994089215822673,
  0.668913398094888, 0.101781714839008, 0.60802422493822, 0.0428021497472084, 
    1.02805127557532, 0.0744361837379512, 0.145260655714142, 
    0.0660277311001161, 0.0908284957784663, 0.092030354084127,
  0.605472357185923, 0.111315582292847, 0.651872679199107, 
    0.0429375119918619, 1.06859706358131, 0.0893670462114645, 
    0.1257249072332, 0.0772872252907215, 0.0888755163010211, 
    0.0821474116371171,
  0.697649773470197, 0.0996571963622462, 0.639252686868213, 
    0.0362943524721688, 1.14405243295968, 0.0749034710578507, 
    0.128102274047438, 0.0754736676904394, 0.0870332345860361, 
    0.0907967628269082,
  0.642842305041659, 0.104780375371438, 0.628323465586934, 
    0.0404525010322863, 1.07903577993298, 0.0728212020820249, 
    0.115237092205659, 0.0527236917377181, 0.0879209397205564, 
    0.0747098676138943,
  0.704165526190996, 0.101149836067291, 0.687332178386382, 
    0.0608049907309955, 1.12040604602414, 0.0774964759079234, 
    0.129761968119214, 0.0485261149361954, 0.0940265066596164, 
    0.0782602771756522,
  0.670391594749706, 0.0856165809975813, 0.65844701276798, 
    0.0485677725572783, 1.0781430965939, 0.067805504685918, 
    0.134669322378191, 0.0616566841756565, 0.0901612451161968, 
    0.0701490703176623,
  0.692825351665683, 0.0990939436317027, 0.584608407666883, 
    0.0464301144944701, 1.10331879528144, 0.0856574801001614, 
    0.120839767874022, 0.0699192061755195, 0.0751823091557432, 
    0.0901252619251056,
  0.744847705592634, 0.0956145276534496, 0.609284245785288, 
    0.049329727451719, 0.997197719430287, 0.073260956918216, 
    0.126229083940129, 0.0696543574363107, 0.0898893015346432, 
    0.0894965744353479,
  0.636273592664875, 0.098951572757285, 0.580173816364282, 
    0.0588743058901234, 1.04155806962804, 0.0624669365377144, 
    0.131802300654908, 0.0684808186590922, 0.0886159931519006, 
    0.0933489791739082,
  0.663360109357266, 0.102976204910454, 0.593206101367186, 
    0.0631187737095126, 1.08656543352393, 0.0808064357219051, 
    0.138927229532029, 0.0640716419443061, 0.0836263270797862, 
    0.105101974204479,
  0.692381357004722, 0.106769355034358, 0.718649477345344, 
    0.0502400805144417, 0.977070920269999, 0.0825064153477936, 
    0.131008855448697, 0.0654173355190461, 0.0835547911374756, 
    0.0824074892346797,
  0.690585545674835, 0.0993092258024292, 0.635608630748956, 
    0.0426362755687328, 1.0187924493771, 0.0644436855117654, 
    0.13152270816941, 0.0629879022684827, 0.0915138659079038, 
    0.0977355475980404,
  0.740224462418991, 0.0903568276268019, 0.640083170458828, 
    0.0531144662615762, 1.02351867934167, 0.0883034669729905, 
    0.121507673772112, 0.0718772328396006, 0.085580944734258, 
    0.0917875107857166,
  0.673455578286775, 0.0965865703930499, 0.711093393205674, 
    0.035560975325555, 1.12511975048084, 0.059860351331803, 
    0.128488680527436, 0.0721128112681947, 0.0826642978509311, 
    0.0900534896563905,
  0.664735476023624, 0.0873380021345173, 0.623132314633577, 
    0.0571430435192994, 1.05015326660781, 0.0918165409717349, 
    0.125844522249483, 0.0530362180528401, 0.0848934332768399, 
    0.0819476988517322,
  0.600242143313784, 0.0886476330872139, 0.552488839879997, 
    0.0259021058285113, 1.0512113593493, 0.0724292994964121, 
    0.124203997748912, 0.059887783331052, 0.0874129592975392, 
    0.0851885532956717,
  0.585295030993011, 0.089453872588872, 0.614764785472634, 
    0.0558694085689731, 1.06661795528085, 0.0928464303703535, 
    0.114777863744957, 0.0688321141807997, 0.0713587888833514, 
    0.0811343365077226,
  0.65912368744219, 0.0996309088654399, 0.641319508329545, 
    0.0615769501157913, 1.08230324551134, 0.0567238985926939, 
    0.136619304830285, 0.0788038786133533, 0.0906581410152499, 
    0.086139503728756,
  0.670094034246549, 0.104412015500271, 0.632701345433991, 
    0.0477881699899856, 1.034912770081, 0.0802794521354041, 
    0.120563826621629, 0.0689717096407206, 0.0849125248803306, 
    0.0917886229301078,
  0.682827757271712, 0.107251195365199, 0.66777437999907, 0.0449484403155853, 
    1.03360471019157, 0.0742721772835777, 0.125591392550819, 
    0.070017352609201, 0.0857285835434776, 0.0858332308424288,
  0.667861533746507, 0.112897791583198, 0.588063400739635, 
    0.0429888116370301, 0.998138566658631, 0.0722543199589607, 
    0.131185648706548, 0.0675076797806691, 0.0729832259484812, 
    0.0999340826522686,
  0.617805082195423, 0.111369717919059, 0.674364232788444, 
    0.0601755411865058, 1.09142051622498, 0.076619584105231, 
    0.131363756571932, 0.0717907774133309, 0.0859106145410863, 
    0.0824073310876204,
  0.579944282258113, 0.0916550337114139, 0.640432110204853, 
    0.0365472253210639, 1.0840897292827, 0.0611224775976067, 
    0.140441659145725, 0.0709342532192875, 0.0808821772241903, 
    0.093581427467525 ;

 source_phase =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 wind =
  18.8878616178245, 20.5105997593991, 18.8643954886542, 20.9501667515465, 
    23.465771443739, 22.087862753995, 17.9456103707668, 19.6882836864023, 
    24.7693145760203, 18.7380529638129,
  23.2522038244511, 20.6111502509785, 20.4311122947025, 23.1308938989109, 
    24.387687822062, 22.2483901167309, 20.617652069705, 20.5089141235035, 
    23.9492298966891, 22.6035276954575,
  18.9240901435263, 22.231258602196, 17.8474406689875, 20.2118053081679, 
    22.7891223577641, 20.67017734292, 19.3233980030139, 21.8862433684642, 
    20.7913777894508, 18.9057007934982,
  19.844746542308, 21.4997188979208, 19.6203138690629, 18.974735253704, 
    22.5572866044105, 22.9696164377175, 21.8336354881495, 21.7164660297489, 
    23.2915228644894, 22.6084196625979,
  20.7432116666115, 18.4459807650847, 19.9446722044031, 20.6203923927682, 
    23.4372276367945, 23.3805321014444, 20.1811367362091, 21.1631742932128, 
    22.1093202313184, 19.9136179586323,
  22.9407036460927, 20.7375580363566, 20.031031558881, 22.2151150595632, 
    26.845544076927, 22.2076891890542, 19.924842885734, 20.1611581769524, 
    21.7502614299495, 22.1688349576853,
  18.7315500873134, 20.0215366448487, 18.0334534036964, 20.0700313862451, 
    23.8385586052104, 25.0830880415971, 18.344501924879, 18.4406004612989, 
    22.6691885982102, 21.2254878822084,
  19.67475807272, 18.4606795121927, 20.7313733394879, 21.7563957499273, 
    20.4956564979568, 20.6405786327907, 19.105504422694, 21.991105323251, 
    22.1861184014487, 21.7532717674772,
  19.7504492540595, 22.3827877720173, 20.4264047486867, 23.115129937219, 
    24.678706612633, 24.3331828237285, 20.6572510355946, 20.4708863923982, 
    24.1851909384539, 22.1286180761312,
  19.4379967472109, 22.2770609645104, 19.3039364565727, 20.3145090162896, 
    23.3742140665709, 23.5205329173619, 19.299428998702, 20.1092611078559, 
    22.7744806265657, 21.8243402793692,
  22.7307472160906, 22.5201878200996, 19.6909891481612, 19.1518275046323, 
    22.5396704862736, 20.9935363979498, 19.7742714860476, 22.092204372929, 
    22.5398862013232, 21.244269921591,
  20.8040527333727, 19.7062591034469, 20.3012427857018, 21.43831956058, 
    25.1011258388991, 22.3601517554615, 18.5844953055333, 18.4521881184239, 
    22.2187973753926, 20.6539925203781,
  21.9250775414466, 22.1964379648958, 21.1894900678812, 21.0219420553002, 
    23.8320737643352, 22.1784421588297, 22.1230248413386, 23.1903955673574, 
    23.0475329611352, 20.9010840544659,
  22.8916114511298, 19.1788798524568, 19.0523903374973, 22.8319551095694, 
    26.0409685435071, 24.0916355141043, 19.6847843159052, 18.9964668414123, 
    20.5466682279677, 22.465973246003,
  23.7458670667284, 20.384650072923, 20.8749331217953, 21.6125292829048, 
    27.2647881324455, 23.5735935754103, 19.6357927385124, 20.5994093957794, 
    22.8638291063095, 22.8618385453535,
  19.755456640864, 20.084549216035, 21.0063647654413, 18.3333804077587, 
    24.0095306341033, 20.0694107151001, 21.0831404734352, 19.7474231116456, 
    22.5247476019059, 21.3052401614598,
  21.5313455740038, 18.6407658588039, 17.0657757613842, 24.1787684340902, 
    22.1354647026159, 23.3145622405713, 21.9649816417515, 20.8430960940291, 
    20.3828777424838, 21.7719834322644,
  18.8670093681884, 21.8630572831257, 20.7764153686908, 18.7087043859129, 
    22.7308715968205, 22.3167838973348, 19.179701805822, 20.6953641234092, 
    22.6533895473616, 21.2617242605664,
  21.1667196600591, 20.477397692895, 22.9321107150729, 21.1490416434017, 
    23.4287421175976, 25.4730540314341, 22.3023173534885, 19.3680210856072, 
    22.2596192542619, 19.5297804077155,
  18.7863014076052, 19.6587974149866, 20.0949760583844, 21.8179836509743, 
    21.84293090537, 20.1226939725781, 17.2150683554386, 19.4301835377285, 
    21.3647469607722, 19.9757912104126,
  20.7270187601401, 19.8174232570581, 17.8658760370612, 19.6807028249001, 
    25.0590900617703, 21.8262883670294, 20.9774819695221, 21.0340771998763, 
    25.4319238891586, 20.2761460088784,
  17.7953900092841, 19.7339800199595, 20.2272580708095, 20.2799958299291, 
    23.9667860320722, 21.3976533233382, 19.2435246770786, 17.5875991848977, 
    22.3514320335223, 20.1381586156734,
  21.7222850335815, 23.6516335908216, 21.801599908578, 20.5752909401679, 
    26.2737603142129, 23.5819428595612, 19.473073714833, 20.733047509717, 
    25.0868113326582, 22.2194172597872,
  21.2360824967397, 19.6366803638275, 16.5694855052028, 19.6166233414677, 
    20.2578684523165, 21.939233106135, 18.7584379666643, 18.9919746155208, 
    21.7679994316744, 19.1923067898648,
  21.4048888845484, 21.4068144428296, 20.4665271530933, 23.1811126267579, 
    23.3809488207113, 23.5737515845015, 19.174858415579, 19.1530346095299, 
    21.4525001734422, 20.2559807569082,
  21.0218651726912, 20.4477845992378, 19.7761560115001, 21.7084688394341, 
    21.6448090673114, 22.6376819730977, 18.1255223695743, 19.6022637130752, 
    20.7739707105217, 19.8287599174694,
  19.9134240254978, 18.517548881749, 18.5628247276894, 20.7256192129135, 
    23.0991009169285, 20.4452100247519, 18.2139464313708, 18.5612176292671, 
    20.8365754038312, 18.7950063987217,
  21.5197497485678, 21.9987399422141, 20.3354565198331, 20.5682711021745, 
    26.1025913738771, 23.4776218723257, 20.3875066708043, 19.6714772682124, 
    22.7640524955675, 23.0809160290828,
  18.4643296694728, 20.1533319412248, 17.2547116580559, 22.2117819629353, 
    24.813551293135, 24.8690742745485, 19.3597151028828, 20.8446081537042, 
    19.7554255412557, 19.3301350971378,
  19.3729242919544, 19.4016119972136, 18.3944254686152, 21.1241323861084, 
    23.9203408937151, 23.8046374779042, 20.7733997944827, 23.3663679637015, 
    23.4216023885655, 20.9866470161893,
  19.8720168690158, 20.2065059549383, 19.5739653472285, 21.1085329919056, 
    22.391010372193, 22.3169174229268, 20.9287800849837, 20.2863265093175, 
    23.9437066238772, 22.296935235681,
  23.3916905053632, 22.2800023676223, 20.4743795152684, 21.6759297344214, 
    24.9877378001156, 24.2652694841964, 22.0183130845317, 21.6905599238225, 
    20.3144431498968, 22.7509128963856,
  19.5097937926345, 17.7352082364713, 17.7046245109348, 18.9145789813742, 
    22.8824630119069, 20.7202433944725, 17.6258603061018, 21.2029153263524, 
    23.4137282334664, 22.1963302232893,
  20.5174457838452, 20.2862142936556, 17.3969665932354, 21.0802386239695, 
    25.0550266432941, 22.679123077703, 19.7309534528068, 21.2397104449681, 
    20.7277422715523, 19.6193614962424,
  18.829741897392, 18.5877781423972, 19.3293464252882, 19.4985675565328, 
    21.8529908025487, 23.7868665047148, 18.5826397231846, 18.2740382428648, 
    19.7280391848824, 19.1049277294864,
  23.4335790789733, 20.9413789961346, 18.9499980706236, 21.6536185179146, 
    22.1710955576571, 21.2541026434068, 19.69373873595, 19.1457445554472, 
    22.4710199032392, 22.6824707974808,
  19.223850958079, 20.4904915867701, 20.716450835281, 22.8482717220375, 
    23.9191152457699, 22.4735647363965, 20.3531129868459, 19.0325499064905, 
    21.2902314155465, 17.3193900382335,
  20.3540428467933, 23.2469312845439, 19.6210584375343, 18.3372583513546, 
    24.3054738317848, 24.299591137249, 19.899985427815, 20.984058848881, 
    23.5124690566524, 20.0418825152151,
  18.6017578188928, 18.5379525177465, 20.6453901811478, 22.5894952932996, 
    23.4488994041509, 22.3808982388218, 22.3037790764205, 21.4269160813809, 
    20.6903984988513, 21.4263725014155,
  20.7896097616709, 20.1021383770624, 19.7874854000958, 23.9507827718466, 
    23.5770165052486, 23.1797032552146, 18.8294460091907, 20.7625816698803, 
    21.0081805322973, 23.2111034445367,
  21.3108859337444, 22.2443510203523, 22.1200243260722, 22.3737673753213, 
    23.526959848853, 22.8520698373318, 20.2012115129689, 19.9211795839965, 
    21.8568111219802, 21.2602377223271,
  21.3377012812665, 20.5913648552058, 20.8446261046859, 18.978822825826, 
    21.9277537020712, 21.561595483018, 19.3973789324587, 19.9594627909544, 
    21.7711875883914, 19.1844457713265,
  19.9947016186541, 22.2126578708498, 19.3034660987393, 20.3172572279985, 
    23.646044198177, 24.9504497636684, 18.6282329191562, 19.2656602748154, 
    20.4992009238158, 20.3711781016258,
  18.7877932233892, 17.6826964278316, 19.5284570994326, 19.4121465276594, 
    20.7114355849927, 22.4502814063694, 18.5222326504203, 21.7478274031874, 
    21.1083531268589, 19.3787987068081,
  19.8080259275271, 20.8457488755231, 19.7543541329113, 22.3314545823551, 
    21.9109139298451, 24.613020955649, 20.8192771966241, 21.5371498771083, 
    20.0575120457023, 21.7125784558468,
  20.7707881856599, 17.5128639696664, 18.3739587662555, 23.35697998771, 
    21.8375468213202, 22.7910706546636, 18.1650749805324, 20.2911815400024, 
    24.2387365465885, 21.7418683632671,
  21.9534565081831, 18.2681244672551, 20.2008460873529, 18.0745915654848, 
    22.4300144651637, 18.6768382670302, 17.9892256633899, 20.656111196466, 
    21.8944155703138, 20.4480049684079,
  19.8904121769397, 20.6475292774392, 20.7793705633924, 21.2842488784893, 
    21.6790003786855, 24.1688443663261, 21.2246231363445, 20.1765549720723, 
    21.4186618120173, 20.1572631294788,
  20.5170292535676, 19.9327766514699, 17.663831265066, 18.3203339100328, 
    22.8755228218978, 21.2744086677694, 17.65597962265, 20.9710401713313, 
    23.3633038529296, 21.2699119386344,
  19.8592343837555, 18.8320644742668, 20.0875806497597, 21.15338503112, 
    23.4223863695157, 21.5164239986627, 18.5893963481967, 18.0570902430335, 
    22.5737309398729, 21.1900483317734,
  20.6704658362762, 21.2488854205595, 18.7663315451817, 19.4916043935036, 
    23.9640256543887, 25.2032754479913, 20.9091652489286, 23.3912741698398, 
    22.2303670352879, 21.3774986479971,
  23.0427801528253, 21.7554867033045, 19.720097123592, 20.9616757217572, 
    23.8133029249937, 22.617786378956, 22.7669569461707, 21.7779045273193, 
    22.6348553410464, 21.3108210499112,
  18.9676115766632, 20.5849578140449, 19.6538834838259, 19.5734126164061, 
    21.2738355795323, 20.8827920334113, 21.3363412233413, 18.8654641189581, 
    21.9687857496241, 20.7461765683046,
  21.0645990350082, 22.414192144478, 18.0047727426321, 20.5477662704291, 
    23.439653692729, 23.4809993667765, 19.460957559075, 17.8703765785006, 
    22.4291299747626, 22.4986390329008,
  19.7902522344808, 17.6693246218612, 17.8139106461161, 20.9767944770421, 
    20.6862663327826, 21.5353195718665, 17.6352843833129, 20.9121153705479, 
    21.6770022074446, 20.7625711695432,
  16.5284232803164, 19.3906054256954, 18.3762056116535, 19.6534284899208, 
    23.1325747900031, 20.5571633486414, 16.9082342833119, 18.8572859962945, 
    21.4055175823849, 17.4140237414064,
  21.6838465377355, 19.0198069965268, 18.6574579466846, 21.2980110554014, 
    22.5448144535281, 21.6959289624296, 20.9496160142242, 20.2986595043004, 
    21.5980678127403, 23.854726786525,
  20.6483803465252, 21.7449650556957, 21.8487716077131, 19.1210379129678, 
    25.8377036786091, 22.6995170450388, 20.909260580497, 19.4329797310917, 
    23.3645715042855, 21.5253523186528,
  21.1868777352735, 20.2000320015986, 21.4542242986346, 22.3055296327978, 
    21.1278374962575, 20.5678419064391, 21.8054912578213, 22.0736284829024, 
    21.6026972730378, 20.109367978749,
  18.423642100131, 19.6606479449028, 15.4283925169503, 19.6267476462958, 
    21.4924268826484, 22.931028518186, 18.0915925533298, 18.8119144153314, 
    20.0647658794792, 19.2723572851612,
  19.1222115275441, 18.6073639022286, 18.967366488319, 20.7060698070771, 
    22.720224055304, 20.8178110188525, 17.5240227555594, 18.907806714628, 
    21.4522040910744, 20.0050463510553,
  17.6970239471897, 21.8857286474179, 19.2399713490441, 22.5901302902431, 
    23.872656297699, 20.2971028495475, 20.3735492575734, 22.4130848815546, 
    19.5685342285705, 21.3328675331751,
  21.2222582429363, 20.9118896174041, 20.788033310137, 23.0196525454963, 
    26.1393904151394, 23.0590430042083, 21.4134090088275, 20.0966012314036, 
    24.4189425368623, 21.7868448899765,
  22.0114998434758, 23.4530589004457, 20.6212885766811, 21.040969712386, 
    21.2196786494058, 22.5504067162339, 20.9506950741401, 20.0857379913981, 
    21.9959281992724, 21.6651797706408,
  20.8197535720609, 21.3632154513741, 20.827553489744, 24.2169879258077, 
    25.466369138722, 20.694731859809, 19.859471303691, 19.922395069373, 
    21.9275669451139, 23.2748885207702,
  21.0222788055568, 19.9087140088049, 16.977468856117, 20.9239834467574, 
    23.3156602890876, 23.0898309311607, 20.1160769839928, 21.5717294115429, 
    20.9187957551354, 19.8501304687968,
  18.5989900118354, 17.0362835103711, 18.9906956596028, 18.0562546655531, 
    21.7934672794287, 22.1539364819667, 17.3660760689521, 19.2821162488501, 
    21.7619667044534, 21.1891563222287,
  22.4528645620421, 21.0869455084233, 20.3628462075834, 21.6990407865034, 
    26.7107485067987, 22.3221919490598, 21.1194211241627, 22.5615695912112, 
    20.9001728433711, 23.5684054148435,
  19.5929891903761, 21.6815064162502, 19.5141823141361, 19.0659013318649, 
    24.5491137187019, 21.4956908180339, 19.0170526589544, 23.2484406049537, 
    22.7456815923275, 20.1237558593041,
  21.0207938238242, 22.7354582708397, 20.4671283982593, 21.0493980127017, 
    24.937870302882, 22.9330832701693, 18.8346938058637, 21.8390949244266, 
    23.4394771842326, 20.4348629740187,
  22.439495672097, 22.2239780608614, 20.3996842406818, 21.4254754910791, 
    24.106737871831, 23.3119504508935, 20.8994998889703, 22.3330259854594, 
    25.3805125133777, 20.7784963045747,
  20.232245436484, 22.0200202240123, 20.6019164348694, 21.057781977944, 
    23.172636302578, 22.3348181788789, 20.7045228585292, 19.9531735879883, 
    23.2800237633514, 23.5421837505942,
  20.4398067080974, 19.4728201051856, 18.8645151763593, 20.0891442489632, 
    24.7948300744381, 23.1911378224939, 20.2501268835173, 21.7607671966821, 
    22.5906462412284, 19.7597644157044,
  20.9523943879368, 18.4824702937178, 18.8983723120338, 20.0991953081211, 
    22.7030969531206, 22.8413271019972, 18.6095637582357, 18.8571955991314, 
    23.1506791966985, 22.2877092345909,
  16.7887262019891, 18.0019591852751, 18.8797432227189, 19.2664227013896, 
    22.3239973543214, 22.47964177237, 18.9294272110294, 18.2736421940564, 
    22.0823787925044, 17.7387410156788,
  20.5299330334108, 20.5398621007894, 18.0392781050728, 20.1767471005062, 
    22.3865301468366, 21.3057294144812, 21.9069568224142, 20.6382918315267, 
    22.8996383953502, 23.4800623410846,
  20.2609031629648, 19.7067403229904, 20.8511071683591, 21.7238847658687, 
    24.0613342193886, 27.0355837888976, 21.8413687235427, 20.746649554369, 
    22.9266861670549, 21.1312640755266,
  17.2992094461665, 20.6030462497745, 19.6843961359695, 18.9370275547855, 
    22.5458655509215, 21.5522069823609, 21.1690053294, 18.7739085406312, 
    21.5027740403596, 20.3155182551213,
  20.5139437114064, 21.8262510693013, 21.7713537017965, 23.2478336151425, 
    26.6875073678778, 25.0745281358079, 20.0272128845192, 20.7023844831634, 
    23.1838820029332, 22.4006274475935,
  18.272571541994, 19.9991822362101, 22.2440388109405, 19.9216074827898, 
    26.0693016587779, 22.5742468820978, 21.2450006513391, 19.7373964708486, 
    21.7854094808213, 21.2048647004853 ;

 concentration_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 mean_source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_phase_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 source_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wind_priorinf_mean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 concentration_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 mean_source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_phase_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 source_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 wind_priorinf_sd =
  0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6 ;

 location = 0, 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9 ;

 time = 41.666666666666667 ;

 advance_to_time = 41.666666666666667 ;
}
