netcdf perfect_input_saw {
dimensions:
	member = 1 ;
	metadatalength = 32 ;
	location = 10 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double concentration(time, member, location) ;
		concentration:long_name = "tracer concentration" ;
		concentration:units = "mass" ;

	double mean_source(time, member, location) ;
		mean_source:long_name = "mean source" ;
		mean_source:units = "mass/timestep" ;

	double source(time, member, location) ;
		source:long_name = "source" ;
		source:units = "mass/timestep" ;

	double source_phase(time, member, location) ;
		source_phase:long_name = "source phase" ;
		source_phase:units = "radians" ;

	double wind(time, member, location) ;
		wind:long_name = "wind" ;
		wind:units = "gridpoints/timestep" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;
		location:axis = "X" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

// global attributes:
		:title = "true state from control" ;
                :version = "$Id: perfect_input_saw.cdl 11441 2017-04-06 22:00:44Z nancy@ucar.edu $" ;
		:description = "Saw tooth pattern for mean source at grid points 1 3 and 5" ;
		:model = "simple_advection" ;
		:destruction_rate = 5.555556e-05 ;
		:history = "same values as in perfect_ics r3014 (circa July 2007)" ;
data:

 MemberMetadata =
  "true state" ;

 concentration =
  4955.56911479461, 4588.67496000528, 5858.36599874513, 4999.69039456505, 
    7448.19165275393, 6288.13835578302, 5324.11858864165, 4534.00933544095, 
    3680.63282566218, 3271.88221046538 ;

 mean_source =
  1, 0.1, 1, 0.1, 1, 0.1, 0.1, 0.1, 0.1, 0.1 ;

 source =
  0.666265198647732, 0.127551533104185, 0.565544571945061, 
    0.0742006468377414, 1.03224698059521, 0.0787975040071264, 
    0.070861950781954, 0.103574720584732, 0.0391374013868522, 0.12572086939668 ;

 source_phase =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 wind =
  21.848170394285, 20.1481610783294, 20.9302183644107, 20.7697938399321, 
    20.6169818006319, 22.3993132701218, 22.0327241481922, 22.2729309428977, 
    23.2970570683049, 21.3608001247452 ;

 location = 0, 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9 ;

 time = 41.666666666666667 ;

}
